module ElectroMagnet(color, out){
    input [0:width]color;
    output [0:width]out;
}

endmodule